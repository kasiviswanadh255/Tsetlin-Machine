module tb(

    );
    reg [783:0] features;
    reg [1567:0] exclude_state_1,exclude_state_2,exclude_state_3,exclude_state_4,exclude_state_5,exclude_state_6,
    exclude_state_7,exclude_state_8,exclude_state_9,exclude_state_10,exclude_state_11,exclude_state_12,
    exclude_state_13,exclude_state_14,exclude_state_15,exclude_state_16,exclude_state_17,exclude_state_18,
    exclude_state_19,exclude_state_20;
    
    wire verdict;

    IM_INFERENCE DUT (features,exclude_state_1,exclude_state_2,exclude_state_3,exclude_state_4,exclude_state_5,exclude_state_6,
                exclude_state_7,exclude_state_8,exclude_state_9,exclude_state_10,exclude_state_11,exclude_state_12,
                exclude_state_13,exclude_state_14,exclude_state_15,exclude_state_16,exclude_state_17,exclude_state_18,
                exclude_state_19,exclude_state_20,verdict);

        initial
        begin
        exclude_state_1=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_2=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_3=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_4=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_5=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_6=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_7=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_8=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_9=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_10=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_11=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_12=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_13=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_14=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_15=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_16=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_17=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_18=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_19=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        exclude_state_20=~{784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,~784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000};
        
            features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011111000000000000000000000011111100000000000000000000011111111100000000000000000111111111110000000000000000011111110111000000000000000011110010001100000000000000011111000000111000000000000011100000000011100000000000001100000000001110000000000001110000000000111000000000000111000000000011100000000000111000000000011100000000000011100000000011100000000000001110000000011100000000000000111000000111100000000000000011110011111100000000000000001111111111100000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//0
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000111111110000000000000000000111111111111110000000000000111000011111111110000000000011100001111111111100000000001100000110000001110000000000110000000000000001000000000011000000000000000110000000001100000000000000011000000000111000000000000001100000000011100000000000000111000000000110000000000000011000000000011100000000000001100000000001110000000000000110000000000011100000000000111000000000000111000000000111000000000000001110000000111000000000000000011111001111100000000000000000111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//0
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000001111111100000000000000000011111111111110000000000000111111111111111110000000000111111111100011111100000000111111110000000011110000000011111110000000001111000000000111110000000000011100000000011110000000000011110000000011110000000000001111000000001111000000000001111000000000111000000000001111000000000011100000000001111100000000001111000000011111100000000000011111101111111100000000000001111111111111000000000000000001111111111000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//0
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000001111110000000000000000000011111111100000000000000000011111111110000000000000000011111111111000000000000000111111111111100000000000000111111111101110000000000000111111101110111000000000000011110000000011100000000000011111000000001110000000000011110000000000111000000000011111000000000111100000000001111000000000111110000000000111100000000111110000000000011100000000111110000000000001111100001111110000000000000111111111111100000000000000011111111111100000000000000000111111111100000000000000000001111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//0
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000111111000000000000000000000111001110000000000000000000111000011000000000000000000111100001100000000000000000111110000011000000000000000111110000001100000000000000011011000000110000000000000011101100000011100000000000001100010000001110000000000000110000000000111000000000000111000000000011000000000000011100000000001100000000000000110000000000110000000000000011000000000110000000000000001100000000111000000000000000111000000111000000000000000001111111111000000000000000000011111111000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//0
        
//        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000011000000000000000000000000011100000000000000000000000001110000011000000000000000000110000001100000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000110000000000000000000000000001110000000000000000000000000011111000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        
//        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000111111111111110000000000000111111111111111100000000000111111111111111110000000000111111111111111111000000000011111111111111111110000000001111111111111111111100000000111111111111111111110000000011111111100000011111000000001111111110000001111100000000111110000000000111110000000011111000000000111111000000001111100000000111111000000000111110000000111111100000000011111000000111111110000000001111100001111111111000000000111111111111111111000000000011111111111111111000000000000111111111111111100000000000001111111111111100000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        

        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000001111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011110000000000000000000000001111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000111100000000000000000000000111100000000000000000000000011100000000000000000000000011110000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000001111000000000000000000000000111100000000000000000000000111100000000000000000000000011110000000000000000000000011110000000000000000000000001111000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001111000000000000000000000000111110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111100000000000000000000000011110000000000000000000000001111000000000000000000000000111110000000000000000000000011111000000000000000000000000111100000000000000000000000011110000000000000000000000000111000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000110000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        
        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000000110000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000111000000000000000000000000011000000000000000000000000001100000000000000000000000000110000000000000000000000000011000000000000000000000000001110000000000000000000000000111000000000000000000000000011100000000000000000000000001110000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        

//        #20 features = 784'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000011100011100000000000000000001110011110000000000000000000111001111000000000000000000011110111000000000000000000001111111100000000000000000000111111100000000000000000000001111100000000000000000000000111110000000000000000000000011110000000000000000000000011111000000000000000000000001111100000000000000000000001111110000000000000000000000111111000000000000000000000111111110000000000000000000011111111000000000000000000011111111100000000000000000001111111110000000000000000000111111111000000000000000000011111111100000000000000000001110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;//1        


        #20 $finish;
    end
endmodule
